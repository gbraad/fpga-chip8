3C
7E
C3
C3
C3
C3
C3
C3
7E
3C
00
00
00
00
00
00
3C
18
18
18
18
18
18
58
38
18
00
00
00
00
00
00
FF
FF
60
30
18
0C
06
C3
7F
3E
00
00
00
00
00
00
3C
7E
C3
03
0E
0E
03
C3
7E
3C
00
00
00
00
00
00
06
06
FF
FF
C6
66
36
1E
0E
06
00
00
00
00
00
00
3C
7E
C3
03
FE
FC
C0
C0
FF
FF
00
00
00
00
00
00
3C
7E
C3
C3
FE
FC
C0
C0
7C
3E
00
00
00
00
00
00
60
60
60
30
18
0C
06
03
FF
FF
00
00
00
00
00
00
3C
7E
C3
C3
7E
7E
C3
C3
7E
3C
00
00
00
00
00
00
7C
3E
03
03
3F
7F
C3
C3
7E
3C
00
00
00
00
00
00
