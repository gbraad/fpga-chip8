	.INIT_08(256'h1636E826E846A2E08268785FEA065FEA1808F033223233267666642242332311),
	.INIT_09(256'h0F21F29266926851F3F2AE063258FC0258FC086FEA7103E2DDBD2A6236060676),
	.INIT_0A(256'hBD2AD1B1F4B104B104180808B8080898D1A1F4A104A104180808A80808882104),
	.INIT_0B(256'h0104180808D808089851E1F4E104E104180808C80808889236E806E8F6BD0676),
	.INIT_0C(256'hA292683103E878E846DDBD2A62C236519216E826E8C6DD3606DD2A5101F40104),
	.INIT_0D(256'hAA6D8A516307076DAA6D8AD103C2066DAA6D8A0606160602EA262602EA1626E0),
	.INIT_0E(256'h6DAA6D8A9103F7F76DAA6D8AD103C2066DAA6D8A7123076DAA6D8AD103C2066D),
	.INIT_0F(256'h0671AE0651AE0641AE069888E80678116DCA6DAA51B103F76DAA6D8AD103C206),
	.INIT_10(256'h4838E8F662F104C104A104E82806A103E80608D25848F7040704F704070481AE),
	.INIT_11(256'h0608D207584821F7060103E80608D2F758482107060103E80608D20758486158),
	.INIT_12(256'h040F06075D3A5F38E8F6E0F89D6221F7060103E80608D2F758482107060103E8),
	.INIT_13(256'h04311F1FF6E836F103E8F6D2D8C8E806E103E8F6D2B8A8075D3A5F38E8F6311F),
	.INIT_14(256'h03E1030F86E0BDF7040704F7040704BD3103E8F62AD2B8A8E806787831060476),
	.INIT_15(256'h039104B898E8B103C104A888E1E8B103C104A888E881039104B89861030808E1),
	.INIT_16(256'hBDE1043826E02806E8F6BDF7BDE1043816E02806E8F6BD07BDE1043846E1E881),
	.INIT_17(256'h06010408BD21E8E806F10318FCE02806E8F6BDF7BDE1043886E02806E8F6BD07),
	.INIT_18(256'h2AD2D8C8E8367878E028E8F6BDF706E1040821070611040821070611040821F7),
	.INIT_19(256'hE8A103C104D89891040808110311030F86E0DDF7140724F7040734DD5103E8F6),
	.INIT_1A(256'hC6E8DD07DD1104384611E8A103C104D898E8E103F104C88811E8E103F104C888),
	.INIT_1B(256'h3886E02826E8C6E8DD07DD11043826E02806E8C6E8DDF7DD11043816E02836E8),
	.INIT_1C(256'h073641040851F796310408DD41E8E836E8210318FCE02816E8C6E8DDF7DD1104),
	.INIT_1D(256'h1FEA0808080704E806988808E80678E028E846DDF7061104085107A641040851),
	.INIT_1E(256'h3D1F4A0808E8D23828063828E08183075F1F1F1F1FEA6F1F1F1F1F8A06E0F89D),
	.INIT_1F(256'hE0F1AE065F086FEAE06F1F1F1FEA08080808080808080707A1E0440728A18307),
	.INIT_20(256'h064104E80458E6180848077D3F01E83828210458262104E8045816180848066F),
	.INIT_21(256'h045806180848077D3F51E838286104E8045866180848077D3F31E83828410458),
	.INIT_22(256'h5FEAE0043818B103E00428086FEAE05FEA0703E86FEAE07D3F077D3F71E83881),
	.INIT_23(256'h370007301365511013776620000000E006E0C1033816C10338D1AE16F606E8E0),
	.INIT_24(256'h0000000000000000767743101155631026677310136773101377731010777210),
	.INIT_25(256'h0008000F8888888F000088880000000F00000088000800000000000000000000),
	.INIT_26(256'h0C0000E00E0000600C0000E00E00006000000000000000000000000000000000),
	.INIT_27(256'h000C003009006090030C00300900600000000000000000000000000000000000),
	.INIT_28(256'h0D0B000060C0B0E00E0B060C0000B07000000000000000000000000000000000),
	.INIT_29(256'h000C00609E30C0B00B0609E30C00600000000000000000000000000000000000),
	.INIT_2A(256'h000900F00B007000000D00B00F0030000D07000000000000000000000000D070),
	.INIT_2B(256'h0D0060000000000000000000000C007000000000000090600C03000000000000),
	.INIT_2C(256'h0000000000000000000000000000000000000090000E00F00F00E00003000000),
	.INIT_2D(256'h000000000000000000000000000000000900B0000003009003009000000B0030),
	.INIT_2E(256'h0F0F0F81080C0C894224A5A52442810030F0F0F08000E010C0E0B0F0E0C010E0),
	.INIT_2F(256'h000000000000000000000000000000000F0F0F81C88C0C89C2E4E5E7E7C38100),
