3C
7E
C3
C3
C3
C3
C3
C3
7E
3C
00
00
00
00
00
00
18
38
58
18
18
18
18
18
18
3C
00
00
00
00
00
00
3E
7F
C3
06
0C
18
30
60
FF
FF
00
00
00
00
00
00
3C
7E
C3
03
0E
0E
03
C3
7E
3C
00
00
00
00
00
00
06
0E
1E
36
66
C6
FF
FF
06
06
00
00
00
00
00
00
FF
FF
C0
C0
FC
FE
03
C3
7E
3C
00
00
00
00
00
00
3E
7C
C0
C0
FC
FE
C3
C3
7E
3C
00
00
00
00
00
00
FF
FF
03
06
0C
18
30
60
60
60
00
00
00
00
00
00
3C
7E
C3
C3
7E
7E
C3
C3
7E
3C
00
00
00
00
00
00
3C
7E
C3
C3
7F
3F
03
03
3E
7C
00
00
00
00
00
00
