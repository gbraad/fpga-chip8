	.INIT_08(256'h04E1163104E11631046FF6E12621F4E11621046FF6F65A11D2D2B2521202F0E0),
	.INIT_09(256'h060606E1267104E12671046F06065F0606BA0000E0E12651F4E1164104E11641),
	.INIT_0A(256'hC1046F3F3AE60000E0E126A104E126A104E1269104E12691046F060606065F06),
	.INIT_0B(256'h060104E106F104088686E106E104E106E1F4087686E0E116D104E116C104E116),
	.INIT_0C(256'h4104E1063104087686E1062104E10621F4188686E1061104E1061104187686E1),
	.INIT_0D(256'h815408F6A6E10671A40806A6E10661A408F6A6E1065104E10651F4088686E106),
	.INIT_0E(256'h08E116B104E116B1240856E116A104E116A1A408E1169104E116915408A6E116),
	.INIT_0F(256'h4D3F074D3F06066F3F3AE0E106E1041DE106E1041D0606E0E116D104E116C114),
	.INIT_10(256'h0000000CCCC8E02183071DE02143071D06762206062236062206063A114D3F07),
