	.INIT_08(256'h22C3D0E211C3C0620053F4C300A2F1C3C0220050F1F08202622342C22284F000),
	.INIT_09(256'h728190C320A201C3102290510100508190023210E0C30062F4C3F0E233C3E062),
	.INIT_0A(256'h4220523054F00000E0C360E263C3506272C340E281C330629053030201005363),
	.INIT_0B(256'h50231FC340A201410100C330C20FC32042F141F100E0C3B04292C3A0C231C390),
	.INIT_0C(256'h431FC3A0C31171F100C390E30FC38063F0501100C370831FC360031050F100C3),
	.INIT_0D(256'h435131F1A0C3F063A111A100C3E083A121F1A0C3D0A30FC3C023F1711100C3B0),
	.INIT_0E(256'h60C360E31FC35063A06050C340A30FC3302380E0C320831FC3100340E0A0C300),
	.INIT_0F(256'hA30193A300A4A3523054E0C310A31F10C300030F101110E0C380030FC3708350),
	.INIT_10(256'h0000000DDDD0E0A4001010E00401111001F0040100A4F100A401004402A30293),
