	.INIT_08(256'h8948177E270E870067363750685051283130F0197D8F81072525750E3000E2A2),
	.INIT_09(256'h70C207484E480E02760710100624F48524F4055068E20E238C8A89274D4C0B0A),
	.INIT_0A(256'h8A8922C2F0C210C200506161016060002202F002100200506161016060002300),
	.INIT_0B(256'hA3005061610160600062E2F0E210E20050616101606000482E174E273E8A0B0A),
	.INIT_0C(256'h48480E42002000370E8C8A892728F062489E170E27FE8C4D4C8C8962A3F0A310),
	.INIT_0D(256'h0B040BA3044544050B040B830E2830050B040BF7160504082807460848474600),
	.INIT_0E(256'h050B040B8304C5C4050B040B830E2830050B040BA3D646050B040B830E283005),
	.INIT_0F(256'h7E441E8EC41E3E441E6E0504233E03A2050B050BA38316C6050B040B830E2830),
	.INIT_10(256'h081727CE27E4724462C45222007E4400208E02070100C4134423C5034533C41E),
	.INIT_11(256'h8E020740010004C5034400208E0207C101000445334400208E02074101002709),
	.INIT_12(256'h0070511684095010200EE00E882704C4134400208E0207C00100044423440020),
	.INIT_13(256'h13645080F0370E6400200E07010037CE4400200E0701004684895010200E6481),
	.INIT_14(256'h046501710EE08ACA424A82CB024BC28A6500200E8907010022CE030264042344),
	.INIT_15(256'h03E50F5303376503E50F530365376503E50F5303376503E50F5303850FE30165),
	.INIT_16(256'h8A65012103E01702273E8ACB8A65012103E017C2273E8A4B8A65012103653765),
	.INIT_17(256'h42460FE08A053237CE65002001E01742273E8ACA8A65012103E01782273E8A4A),
	.INIT_18(256'h89070100220E0302E017273E8ACB02E50FE0664A82C60FE0664BC2060FE066CA),
	.INIT_19(256'h37E603860F5303060FE30167046701710EE08CCC024C02CD024D028CE600200E),
	.INIT_1A(256'hFE378C4D8C670121036737E603860F5303372603C60F530367372603C60F5303),
	.INIT_1B(256'h2103E0170227FE378C4C8C67012103E0170227FE378CCD8C67012103E0170227),
	.INIT_1C(256'h4D02270FE087CC02670FE08C8632370E3787002001E0170227FE378CCC8C6701),
	.INIT_1D(256'hE088E0E0E01001214E4101E0203E00E01727FE8CCD02E70FE0874C02E70FE087),
	.INIT_1E(256'h42E009E0E020470100FE3332E0870E1E53EEEEEEEE0B53EEEEEEEE090EE00E88),
	.INIT_1F(256'hE0A7101050605068E050E0E1E10BE1E1E1E1616160604140E7E0034332E70242),
	.INIT_20(256'h35E80F520F5385030234C6A604A8440100680F5275680F520F53050302341E51),
	.INIT_21(256'h0F53A5030234C6A604A8440100E80F520F5345030234C6A60428440100E80F52),
	.INIT_22(256'h5148E00F5E0EC80EE00F5E0E5328E05128100F415128E0A601C6A604A8440188),
	.INIT_23(256'hCEF7FEC0CEFDDEC0CEF73320050000E01EE0A8004001A80141E81201F3F23EE0),
	.INIT_24(256'h0088000000080000F3F79EC0CEDDFEC02337FEC0C0FFF2C0EF808FE0C6BFF6C0),
	.INIT_25(256'h0000000000000000000000000000000000000000000000000000000000000000),
	.INIT_26(256'hA55555555555555AA55555555555555AD88888888888888CD88888888888888C),
	.INIT_27(256'hA5A5655AA5555A5555A5555AA5565A5AA5D8885DC5F88C5FE5D8885DC5F88C5A),
	.INIT_28(256'hA55555555A555555555555A55555555AA5F5F8888C885F888885F8C888885F5A),
	.INIT_29(256'hF5F5555A555A55555055A555A5555F5FA5D8888C5F5D885F85F8C5F5D8888C5A),
	.INIT_2A(256'hA5A5555555555F8CD885555555555A5A7455F85F85F85D8888C5F85FE5F85547),
	.INIT_2B(256'hA5565A5F8888885F85F8888885A5655AA5F88C5D888C555AA555D888C5D8885A),
	.INIT_2C(256'hA5F85F888885DC5F85DC5F888885F85AA5DC5A55555555555555555555A5DC5A),
	.INIT_2D(256'hF888888888888F88888F888888888888A55555555555AA5555AA55555555555A),
	.INIT_2E(256'h080E0F0F03000F00060F0D0F0F06000FF0F0F1033170713294594B4B49840201),
	.INIT_2F(256'h00000000000000000000000000000000080E0F0F03000F0000070F0F0F0F0F0F),
