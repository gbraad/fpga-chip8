F0
90
90
90
F0
00
00
00
70
20
20
60
20
00
00
00
F0
80
F0
10
F0
00
00
00
F0
10
F0
10
F0
00
00
00
10
10
F0
90
90
00
00
00
F0
10
F0
80
F0
00
00
00
F0
90
F0
80
F0
00
00
00
40
40
20
10
F0
00
00
00
F0
90
F0
90
F0
00
00
00
F0
10
F0
90
F0
00
00
00
90
90
F0
90
F0
00
00
00
E0
90
E0
90
E0
00
00
00
F0
80
80
80
F0
00
00
00
E0
90
90
90
E0
00
00
00
F0
80
F0
80
F0
00
00
00
80
80
F0
80
F0
00
00
00
