18
3C
66
C3
FF
C3
C3
C3
C3
C3
00
00
00
00
00
00
FC
FE
C7
C3
FE
C7
C3
C3
FF
FE
00
00
00
00
00
00
3E
7F
E1
C0
C0
C0
C0
C1
FF
7E
00
00
00
00
00
00
FC
FE
C7
C3
C3
C3
C3
C3
FF
FE
00
00
00
00
00
00
FF
FE
C0
C0
F8
C0
C0
C1
FF
FF
00
00
00
00
00
00
FF
FE
C0
C0
F8
C0
C0
C0
C0
C0
00
00
00
00
00
00
